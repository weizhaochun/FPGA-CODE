module dazuoye( clk,led0,led1,led2,rst,en,two);input clk,rst,en,two;output [2:0]led0;output [2:0]led1;output [1:0]led2; reg [2:0]led0;reg [2:0]led1;reg [1:0]led2;reg [31:0]count;reg  clk1;reg[3:0]q=4'b0000;reg[3:0]s=4'b0000;reg[1:0]r=2'b00;always@(posedge clk)begin if(count<=12999999)  count<=count+1;  else  begin  count<=0;clk1<=~clk1;end end    always@(posedge clk1 )if(rst) begin q<=0;s<=0;r<=0;endelse if(en)begin  q<=q;s<=s;r<=r;endelse if(q<=7)   q<=q+1;   else    begin   	 q<=0;	    if(s<=5)	      s<=(!two)?s+1:s;		 else		    begin		     s<=0;			  if(r<=3)			    r<=r+1;			  else			     r<=0;			 end	 end	   always@(q) case(q) 4'b0000:led0<=3'b000; 4'b0001:led0<=3'b001; 4'b0010:led0<=3'b010; 4'b0011:led0<=3'b011; 4'b0100:led0<=3'b100; 4'b0101:led0<=3'b101; 4'b0110:led0<=3'b110; 4'b0111:led0<=3'b111; default:led0<=3'b000; endcasealways@(s) case(s) 4'b0000:led1<=3'b000; 4'b0001:led1<=3'b001; 4'b0010:led1<=3'b010; 4'b0011:led1<=3'b011; 4'b0100:led1<=3'b100; 4'b0101:led1<=3'b101; default:led1<=3'b000; endcasealways@(r) case(r) 2'b00:led2<=2'b00; 2'b01:led2<=2'b01; 2'b10:led2<=2'b10; 2'b11:led2<=2'b11; endcaseendmodule 